#timeunit 1ns
#timeprecision 1ps


module col #(
)
   (
   )
endmodule

